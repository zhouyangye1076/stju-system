`include"conv_struct.vh"
module Multiplier #(
    parameter LEN = 32
) (
    input clk,
    input rst,
    input [LEN-1:0] multiplicand,
    input [LEN-1:0] multiplier,
    input start,
    
    output [LEN*2-1:0] product,
    output finish
);

    localparam PRODUCT_LEN = LEN*2;
    logic [LEN-1:0] multiplicand_reg;
    logic [PRODUCT_LEN-1:0] product_reg;

    localparam CNT_LEN = $clog2(LEN);
    localparam CNT_NUM = LEN - 1;
    typedef enum logic [1:0] {IDLE, WORK, FINAL} fsm_state;
    fsm_state fsm_state_reg;
    logic [CNT_LEN-1:0] work_cnt;

    logic [LEN-2:0] low_product_result;
    logic [LEN:0] high_product_result;
    
    // fill the code
    
endmodule
`ifndef __BUS_STRUCT__
`define __BUS_STRUCT__

package BusPack;

    typedef enum logic [1:0] {OKAY, EXOKAY, SLVERR, DECERR} resp_t;

endpackage

`endif
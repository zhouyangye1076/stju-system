`ifdef VERILATE
    localparam FILE_PATH = "testcase.hex";
`else
    localparam FILE_PATH = "D:\\txt\\system2\\sys-project\\src\\project\\build\\verilate\\testcase.hex";
`endif
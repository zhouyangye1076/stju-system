`ifdef VERILATE
    localparam DATA_FILE_PATH = "initial_data.hex";
`else
    localparam DATA_FILE_PATH = "D:\\txt\\system2\\sys1-sp24\\repo\\sys-project\\lab4-1\\syn\\initial_data.hex";
`endif
`ifdef VERILATE
    localparam FILE_PATH = "testcase.hex";
`else
    localparam FILE_PATH = ;
`endif